module top();












endmodule
