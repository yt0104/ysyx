`define     ISA_WIDTH       64
`define     REG_ADDR_WIDTH  5
`define     AXI_enable 

parameter inst_ecall = 12'd1;
parameter inst_mret = 12'd2;

