`define     ISA_WIDTH       64
`define     REG_ADDR_WIDTH  5
`define     IDUf_WIDTH      7



parameter inst_ecall = 12'd1;
parameter inst_mret = 12'd2;


//`define     ICACHE_enable
//`define     DCACHE_enable







