//负责根据控制信号对数据进行执行操作, 并将执行结果写回寄存器或存储器
module EXU();


endmodule